-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
-- CREATED		"Tue Oct 18 09:21:45 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Block1 IS 
	PORT
	(
		CLK_50M :  IN  STD_LOGIC;
		continu :  IN  STD_LOGIC;
		start_stop :  IN  STD_LOGIC;
		in_freq_anemometre :  IN  STD_LOGIC;
		raz_n :  IN  STD_LOGIC;
		data_valid :  OUT  STD_LOGIC;
		data_anemometre :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END Block1;

ARCHITECTURE bdf_type OF Block1 IS 

COMPONENT counter
	PORT(in_freq : IN STD_LOGIC;
		 raz_n : IN STD_LOGIC;
		 counter : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT diviseur
	PORT(clk : IN STD_LOGIC;
		 clk_1hz : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT mode_fonctionnement
	PORT(clk : IN STD_LOGIC;
		 continu : IN STD_LOGIC;
		 start_stop : IN STD_LOGIC;
		 internal_reset : IN STD_LOGIC;
		 data_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data_valid : OUT STD_LOGIC;
		 data_anemometre : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT edge_detector
	PORT(clk : IN STD_LOGIC;
		 f_in : IN STD_LOGIC;
		 edge : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;


BEGIN 



b2v_inst : counter
PORT MAP(in_freq => in_freq_anemometre,
		 raz_n => raz_n,
		 counter => SYNTHESIZED_WIRE_1);


b2v_inst2 : diviseur
PORT MAP(clk => CLK_50M,
		 clk_1hz => SYNTHESIZED_WIRE_2);


b2v_inst4 : mode_fonctionnement
PORT MAP(clk => CLK_50M,
		 continu => continu,
		 start_stop => start_stop,
		 internal_reset => SYNTHESIZED_WIRE_0,
		 data_in => SYNTHESIZED_WIRE_1,
		 data_valid => data_valid,
		 data_anemometre => data_anemometre);


b2v_inst6 : edge_detector
PORT MAP(clk => CLK_50M,
		 f_in => SYNTHESIZED_WIRE_2,
		 edge => SYNTHESIZED_WIRE_0);


END bdf_type;